// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition"
// CREATED		"Sat Aug 27 16:25:10 2022"

module SEU_ROY(
	ref_clock,
	pll_out,
	out
);


input wire	ref_clock;
input wire	pll_out;
output wire	[7:0] out;

wire	SYNTHESIZED_WIRE_0;





counter	b2v_inst(
	.reset(ref_clock),
	.clk(SYNTHESIZED_WIRE_0),
	.out(out));

assign	SYNTHESIZED_WIRE_0 = ref_clock & pll_out;


endmodule
